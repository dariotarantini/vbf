module main

struct Instruction {
mut:
    operator int
	operand int
}
